`timescale 1ns/1ns
`include"q2.v"
module q2_tb;
reg a,b,c,d;
wire k1,k2,k3,k4;
q2 uut(a,b,c,d,k1,k2,k3,k4);
initial begin
$dumpfile("q2_tb.vcd");
$dumpvars(0,q2_tb);

a=0;
b=0;
c=0;
d=0;
#20;

a=0;	
b=0;
c=0;
d=1;
#20;

a=0;
b=0;
c=1;
d=0;
#20;

a=0;
b=1;
c=0;
d=0;
#20;

a=0;
b=0;
c=1;
d=1;
#20;

a=0;
b=1;
c=0;
d=1;
#20;

a=0;
b=1;
c=1;
d=0;
#20;

a=0;
b=1;
c=1;
d=1;
#20;

a=1;
b=0;
c=0;
d=0;
#20;

a=1;
b=0;
c=0;
d=1;
#20;

a=1;
b=0;
c=1;
d=0;
#20;

a=1;
b=0;
c=1;
d=1;
#20;


a=1;
b=1;
c=0;
d=0;
#20;

a=1;
b=1;
c=0;
d=1;
#20;

a=1;
b=1;
c=1;
d=0;
#20;

a=1;
b=1;
c=1;
d=1;
#20;

$display("test complete");
end
endmodule
	

