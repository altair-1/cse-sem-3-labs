`timescale 1ns/1ns
`include"q3.v"
module q3_tb;
reg a,b,c,d;
wire f;
q3 uut(a,b,c,d,f);
initial begin
$dumpfile("q3_tb.vcd");
$dumpvars(0,q3_tb);

a=0;
b=0;
c=0;
d=0;
#20;

a=0;	
b=0;
c=0;
d=1;
#20;

a=0;
b=0;
c=1;
d=0;
#20;



a=0;
b=1;
c=0;
d=0;
#20;

a=1;
b=0;
c=0;
d=0;
#20;

a=1;
b=0;
c=0;
d=1;
#20;

a=1;
b=0;
c=1;
d=1;
#20;

a=1;
b=1;
c=0;
d=0;
#20;

a=1;
b=1;
c=0;
d=1;
#20;

a=1;
b=1;
c=1;
d=0;
#20;

a=1;
b=0;
c=1;
d=1;
#20;

a=0;
b=1;
c=1;
d=1;
#20;


$display("test complete");
end
endmodule
	

